module imem(
    input [31:0] A,
    output [31:0] RD
);
reg [31:0] RAM [1023:0];

// initial
// $readmemh("riscvtest.txt",RAM);
initial begin
    RAM[0] = 32'h0062E233; //or  x4, x5, x6
    //add x1, x2, x3
    RAM[1] = 32'b0000000_00011_00010_000_00001_0110011; 
    //sub x8, x9, x10
    RAM[2] = 32'b0100000_01010_01001_000_01000_0110011; 
    // and x5, x3, x4
    RAM[3] = 32'h0041F2B3;
    // slt x4, x3, x4
    RAM[4] = 32'h0041A233;  //x4 = (12 < 7) = 0
    //addi x2,x0,5
    RAM[5] = 32'h00500113; //x2 = 5
    //addi x7,x3,-9
    RAM[6] = 32'hFF718393; // x7 = (12 - 9) = 3
    //addi x2,x0,4
    RAM[5] = 32'h00400113; //x2 = 4
    // lw x4, 4(x2)
    RAM[7] = 32'b000000000100_00010_010_00100_0000011; 
    // sw x3, 4(x2)
    //RAM[8] = 32'b0000000_00011_00010_010_00001_0100011; 
    // sw  x6, 8(x9)
    RAM[8] = 32'b0000000_00110_01001_010_01000_0100011;
    //beq x4, x4, 20 
    //RAM[9] = 32'b0000000_00100_00100_000_10100_1100011;
    RAM[9] = 32'h00420A63;
    //add x1, x2, x3
    RAM[10] = 32'b0000000_00011_00010_000_00001_0110011;
    //or  x4, x5, x6
    RAM[11] = 32'h0062E233; 
    //add x1, x2, x3
    RAM[12] = 32'b0000000_00011_00010_000_00001_0110011;
    //or  x4, x5, x6
    RAM[13] = 32'h0062E233; 
    //add x1, x2, x3
    // RAM[14] = 32'b0000000_00011_00010_000_00001_0110011;
    RAM[14] = 32'h3100B3;

end
assign RD = RAM[A[31:2]];

endmodule