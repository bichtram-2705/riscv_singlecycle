module riscvsingle(
    input clk,
    input rst_n,
    output [31:0] PC,
    input [31:0] Instr,
    output MemWrite,
    output [31:0] DataAdr, WriteData,
    input [31:0] ReadData
);

wire [31:0] ALUResult;
wire Zero;

wire PCSrc;
wire [1:0] ResultSrc;
wire [2:0] ALUControl;
wire ALUSrc;
wire [1:0] ImmSrc;
wire RegWrite;

controller controller_ints(
    .Zero(Zero),
    .PCSrc(PCSrc),
    .ResultSrc(ResultSrc),
    .MemWrite(MemWrite),
    .ALUControl(ALUControl),
    .ALUSrc(ALUSrc),
    .ImmSrc(ImmSrc),
    .RegWrite(RegWrite),
    .op(Instr[6:0]),
    .funct3(Instr[14:12]),
    .funct7b5(Instr[30])
);

datapath datapath_ints(
    .clk(clk),
    .rst_n(rst_n),
    .PC(PC),
    .Instr(Instr),
    .ALUResult(DataAdr),
    .WriteData(WriteData),
    .ReadData(ReadData),
    .RegWrite(RegWrite),
    .ImmSrc(ImmSrc),
    .ALUSrc(ALUSrc),
    .ALUControl(ALUControl),
    .ResultSrc(ResultSrc),
    .PCSrc(PCSrc),
    .Zero(Zero)
);
endmodule